
//operation num
localparam NONE = 6'd0;
localparam ADDI = 6'd1;
localparam SLTI = 6'd2;
localparam SLTIU = 6'd3;
localparam ANDI = 6'd4;
localparam ORI = 6'd5;
localparam XORI = 6'd6;
localparam SLLI = 6'd7;
localparam SRLI = 6'd8;
localparam SRAI = 6'd9;
localparam LUI = 6'd10;
localparam AUIPC = 6'd11;
localparam ADD = 6'd12;
localparam SLT = 6'd13;
localparam SLTU = 6'd14;
localparam AND = 6'd15;
localparam OR = 6'd16;
localparam XOR = 6'd17;
localparam SLL = 6'd18;
localparam SRL = 6'd19;
localparam SUB = 6'd20;
localparam SRA = 6'd21;
localparam JAL = 6'd22;
localparam JALR = 6'd23;
localparam BEQ = 6'd24;
localparam BNE = 6'd25;
localparam BLT = 6'd26;
localparam BLTU = 6'd27;
localparam BGE = 6'd28;
localparam BGEU = 6'd29;
localparam LB = 6'd30;
localparam LH = 6'd31;
localparam LW = 6'd32;
localparam LBU = 6'd33;
localparam LHU = 6'd34;
localparam SB = 6'd35;
localparam SH = 6'd36;
localparam SW = 6'd37;
localparam MISC_MEM = 6'd38;
localparam ECALL = 6'd39;
localparam EBREAK = 6'd40;