module invert
(
    input input1,
    output output1
);

    assign output1 = ~input1;

endmodule
